import uvm_pkg::*;
import tests_pkg::*;

module top;

initial begin
    run_test();
end

endmodule